
module mymodule();
    parameter real fc=10e6;
    parameter real bw=25e3;
    analog begin
	// contents of module here
    end
    endmodule
